// list of operations supported by ALU

package operationList;
	const reg[2:0] addop = 0;
	const reg[2:0] subop = 1;
	const reg[2:0] andop = 2;
	const reg[2:0] xorop = 3;
	const reg[2:0] sraop = 4;
	const reg[2:0] load = 5;
	const reg[2:0] store = 6;
endpackage