module ReservationStation(
	input clk,
	output reg[7:0] new_reservationTable[63:0] 
);
	
	
	
	
endmodule