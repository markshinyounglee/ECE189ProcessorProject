// list of operations supported by ALU

package operationList;
	const reg[3:0] add = 4'b0;
	const reg[3:0] sub = 4'b1;
	const reg[3:0] andop = 4'b2;
	const reg[3:0] orop = 4'b3;
	const reg[3:0] load = 4'b4;
	const reg[3:0] store = 4'b5;
endpackage