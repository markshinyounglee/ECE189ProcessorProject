// R-type, I-type, and Memory instructions (LW, SW)

package instructionList;
	typedef rtype[6:0] = 7'b0110011;
	typedef itype[6:0] = 7'b0010011;
	typedef lw[6:0] = 7'b0000011;
	typedef sw[6:0] = 7'b0100011;
endpackage