// R-type, I-type, and Memory instructions (LW, SW)

package instructionList;
	const reg[6:0] rtype = 7'b0110011;
	const reg[6:0] itype = 7'b0010011;
	const reg[6:0] lw = 7'b0000011;
	const reg[6:0] sw = 7'b0100011;
endpackage